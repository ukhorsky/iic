library IEEE;
use IEEE.STD_LOGIC_1164.all;

package parameters is

    constant clk_f : natural := 50; -- MHz
    -- constant iic_scl_
end parameters;

package body parameters is

end parameters;
